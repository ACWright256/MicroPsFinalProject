
//**********************************************************************************************************************************************************//
//																	SPI and MEMORY SECTION																	//
//**********************************************************************************************************************************************************//


//////////////////////////////////////////////////////////////////////
//							SPIWriteMem MODULE						//
//	Contains both the SPI hardware and EBR memory control stuff		//
//////////////////////////////////////////////////////////////////////
/*module SPIWriteMemTest (input  logic clk,
						input  logic sck, 
						input  logic sdi,
						input  logic CE,
						input logic reset,
						input logic get_buffer,
						input logic [5:0] row_0_sel,
						input logic [5:0] row_1_sel,
						output logic sdo,
						output logic [63:0] row_0,
						output logic [63:0] row_1);
	
	
	logic [383:0] data_frame_unpacked;
	logic w_en;
	logic r_en;
	logic [5:0] y_in [63:0];
	
	//get the SPI data into matrix(wire) form
	
	WireArrayToMatrix MatrixStuff(data_frame_unpacked, y_in);
	SPIIn TestSPI(clk, sck, sdi, CE, reset, sdo, data_frame_unpacked, w_en );
	EBRController TestEBR(clk, reset, w_en,r_en,get_buffer, y_in, row_0_sel, row_1_sel, row_0, row_1  );


endmodule*/





//**********************************************************************************************************************************************************//
//																	DISPLAY CONTROL SECTION																	//
//**********************************************************************************************************************************************************//




//////////////////////////////////////////////////////////////////////
//						DISPLAYCONTROLCOLORINPUT	MODULE			//
//							A TESTING MODULE						//
//	Takes in two rows of color data	and drives the display			//
//////////////////////////////////////////////////////////////////////
/*module DisplayControllerColorInput #(WIDTH=4)(input logic clk,
												input logic reset,
												input logic [WIDTH-1:0] r0_map_cm [63:0],
												input logic [WIDTH-1:0] r1_map_cm [63:0],
												input logic [WIDTH-1:0] g0_map_cm [63:0],
												input logic [WIDTH-1:0] g1_map_cm [63:0],
												input logic [WIDTH-1:0] b0_map_cm [63:0],
												input logic [WIDTH-1:0] b1_map_cm [63:0],
												output logic [4:0] current_addr,
												output logic blank,
												output logic latch,
												output logic r0_out,
												output logic r1_out,
												output logic g0_out,
												output logic g1_out,
												output logic b0_out,
												output logic b1_out,
												output logic out_clk,
												output logic read_en);
	//colshift
	logic pwm_en;
	logic [63:0] r0_cm_cs, r1_cm_cs,g0_cm_cs, g1_cm_cs, b0_cm_cs, b1_cm_cs;			
	logic col_cnt_overflow;	
	logic col_sck;
	logic col_cnt_en;	
	//combcolormod
    logic [WIDTH-1:0] pwm_cnt;
	//maprgb
	logic[5:0] ro1_0_sel;
	logic[5:0] ro1_1_sel;
	//ColorModFSM
	logic [4:0] next_addr;
	logic pwm_overflow;
	//////// MainDisplayFSM	////////
	MainDisplayFSM MainDisplayFSMModule(clk, reset, pwm_overflow,current_addr, pwm_en, next_addr,read_en);
	//////// ColorModFSM	////////
	ColorModFSM #(.WIDTH(WIDTH)) ColorModFSMModule(clk, reset, col_cnt_overflow, pwm_en, next_addr,col_sck, blank, pwm_cnt, latch, current_addr, ro1_0_sel, ro1_1_sel, pwm_overflow,out_clk,col_cnt_en);
	//////// CombColorMod	////////
	CombColorMod #(.WIDTH(WIDTH)) CombColorModulationModule(pwm_cnt, r0_map_cm, r1_map_cm, g0_map_cm, g1_map_cm, b0_map_cm, b1_map_cm, r0_cm_cs, r1_cm_cs, g0_cm_cs, g1_cm_cs, b0_cm_cs, b1_cm_cs);
	//////// ColShift	////////
	ColShift ColShiftModule (clk, reset, col_cnt_en,r0_cm_cs, r1_cm_cs, g0_cm_cs, g1_cm_cs, b0_cm_cs, b1_cm_cs, r0_out, r1_out, g0_out, g1_out, b0_out, b1_out, col_cnt_overflow,col_sck);
	
endmodule*/




//////////////////////////////////////////////////////////////////////
//							MemReadDisplay	MODULE					//
//							A TESTING MODULE						//
//////////////////////////////////////////////////////////////////////
module MemReadDisplay #(WIDTH=4)(   input logic clk,
									input logic reset,
									output logic r0_out,
									output logic r1_out,
									output logic g0_out,
									output logic g1_out,
									output logic b0_out,
									output logic b1_out,  
									output logic latch,
									output logic OE,
									output logic sck,
									output logic [4:0] addr);
	
	 
	  logic [63:0] write_buffer [63:0];
	 
	 
	  /*assign write_buffer[0] =  64'b0000000000000000000111111111111111100000000000000000000000000000;
	  assign write_buffer[1] =  64'b0000000000000011111000000000000000011111000000000000000000000000;
	  assign write_buffer[2] =  64'b0000000000001100000000000000000000000000110000000000000000000000;
	  assign write_buffer[3] =  64'b0000000000110000000000000000000000000000001100000000000000000000;
	  assign write_buffer[4] =  64'b0000000001000000000000000000000000000000000010000000000000000000;
	  assign write_buffer[5] =  64'b0000000001000000001110000000000000011100000010000000000000000000;
	  assign write_buffer[6] =  64'b0000000001000000001110000000000000011100000010000000000000000000;
	  assign write_buffer[7] =  64'b0000000001000000000000000000000000000000000010000000000000000000;
	  assign write_buffer[8] =  64'b0000000001000000000000000000000000000000000010000000000000000000;
	  assign write_buffer[9] =  64'b0000000001000000000000111111111110000000000010000000000000000000;
	  assign write_buffer[10] = 64'b0000000001000000000011000000000001100000000010000000000000000000;
	  assign write_buffer[11] = 64'b0000000000100000000011000000000001100000000100000000000000000000;
	  assign write_buffer[12] = 64'b0000000000011000000000111111111110000000011000000000000000000000;
	  assign write_buffer[13] = 64'b0000000000000110000000000000000000000001100000000000000000000000;
	  assign write_buffer[14] = 64'b0000000000000001111100000000000000111110000000000000000000000000;
	  assign write_buffer[15] = 64'b0000000000000000000011111111111111000000000000000000000000000000;
	  assign write_buffer[16] = 64'b0000000000000000000000000011000000000000000000000000000000000000;
	  assign write_buffer[17] = 64'b0000000000000000000000000011000000000000000000000000000000000000;
	  assign write_buffer[18] = 64'b0000000000000000000000000011000000000000000000000000000000000000;
	  assign write_buffer[19] = 64'b0000000000000011111111111111111111111111110000000000000000000000;
	  assign write_buffer[20] = 64'b0000000000000000000000000011000000000000000000000000000000000000;
	  assign write_buffer[21] = 64'b0000000000000000000000000011000000000000000000000000000000000000;
	  assign write_buffer[22] = 64'b0000000000000000000000000011000000000000000000000000000000000000;
	  assign write_buffer[23] = 64'b0000000000000000000000000011000000000000000000000000000000000000;
	  assign write_buffer[24] = 64'b0000000000000000000000000011000000000000000000000000000000000000;
	  assign write_buffer[25] = 64'b0000000000000000000000000011000000000000000000000000000000000000;
	  assign write_buffer[26] = 64'b0000000000000000000000000011000000000000000000000000000000000000;
	  assign write_buffer[27] = 64'b0000000000000000000000000011000000000000000000000000000000000000;
	  assign write_buffer[28] = 64'b0000000000000000000000001100110000000000000000000000000000000000;
	  assign write_buffer[29] = 64'b0000000000000000000000110000001100000000000000000000000000000000;
	  assign write_buffer[30] = 64'b0000000000000000000011000000000011000000000000000000000000000000;
	  assign write_buffer[31] = 64'b0000000000000000001100000000000000110000000000000000000000000000;
	  assign write_buffer[32] = 64'b0000000000000000001100000000000000110000000000000000000000000000;
	  assign write_buffer[33] = 64'b0000000000000000001100000000000000110000000000000000000000000000;
	  assign write_buffer[34] = 64'b0000000000000000001100000000000000110000000000000000000000000000;
	  assign write_buffer[35] = 64'b0000000000000000001100000000000000110000000000000000000000000000;
	  assign write_buffer[36] = 64'b0000000000000000001100000000000000110000000000000000000000000000;
	  assign write_buffer[37] = 64'b0000000000000000001100000000000000110000000000000000000000000000;
	  assign write_buffer[38] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[39] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[40] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[41] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[42] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[43] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[44] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[45] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[46] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[47] = 64'b0000000000000001111000000000000000000000011110000000000000000000;
	  assign write_buffer[48] = 64'b0000000000000001111000000000000000000000011110000000000000000000;
	  assign write_buffer[49] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[50] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[51] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[52] = 64'b0000000000000110000000000000000000000000000011000000000000000000;
	  assign write_buffer[53] = 64'b0000000000000110000000000000000000000000000011000000000000000000;
	  assign write_buffer[54] = 64'b0000000000000110000000000000000000000000000011000000000000000000;
	  assign write_buffer[55] = 64'b0000000000000001100000000000000000000000001100000000000000000000;
	  assign write_buffer[56] = 64'b0000000000000000011000000000000000000000110000000000000000000000;
	  assign write_buffer[57] = 64'b0000000000000000000111111111111111111111000000000000000000000000;
	  assign write_buffer[58] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[59] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[60] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[61] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[62] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[63] = 64'b0000000000000000000000000000000000000000000000000000000000000000;*/


	  assign write_buffer[0] =  64'b1000000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[1] =  64'b1100000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[2] =  64'b1110000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[3] =  64'b1111000000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[4] =  64'b1111100000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[5] =  64'b1111110000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[6] =  64'b1111111000000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[7] =  64'b1111111100000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[8] =  64'b1111111110000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[9] =  64'b1111111111000000000000000000000000000000000000000000000000000000;
	  assign write_buffer[10] = 64'b1111111111100000000000000000000000000000000000000000000000000000;
	  assign write_buffer[11] = 64'b1111111111110000000000000000000000000000000000000000000000000000;
	  assign write_buffer[12] = 64'b1111111111111000000000000000000000000000000000000000000000000000;
	  assign write_buffer[13] = 64'b1111111111111100000000000000000000000000000000000000000000000000;
	  assign write_buffer[14] = 64'b1111111111111110000000000000000000000000000000000000000000000000;
	  assign write_buffer[15] = 64'b1111111111111111000000000000000000000000000000000000000000000000;
	  assign write_buffer[16] = 64'b1111111111111111100000000000000000000000000000000000000000000000;
	  assign write_buffer[17] = 64'b1111111111111111110000000000000000000000000000000000000000000000;
	  assign write_buffer[18] = 64'b1111111111111111111000000000000000000000000000000000000000000000;
	  assign write_buffer[19] = 64'b1111111111111111111100000000000000000000000000000000000000000000;
	  assign write_buffer[20] = 64'b1111111111111111111110000000000000000000000000000000000000000000;
	  assign write_buffer[21] = 64'b1111111111111111111111000000000000000000000000000000000000000000;
	  assign write_buffer[22] = 64'b1111111111111111111111100000000000000000000000000000000000000000;
	  assign write_buffer[23] = 64'b1111111111111111111111110000000000000000000000000000000000000000;
	  assign write_buffer[24] = 64'b1111111111111111111111111000000000000000000000000000000000000000;
	  assign write_buffer[25] = 64'b1111111111111111111111111100000000000000000000000000000000000000;
	  assign write_buffer[26] = 64'b1111111111111111111111111110000000000000000000000000000000000000;
	  assign write_buffer[27] = 64'b1111111111111111111111111111000000000000000000000000000000000000;
	  assign write_buffer[28] = 64'b1111111111111111111111111111100000000000000000000000000000000000;
	  assign write_buffer[29] = 64'b1111111111111111111111111111110000000000000000000000000000000000;
	  assign write_buffer[30] = 64'b1111111111111111111111111111111000000000000000000000000000000000;
	  assign write_buffer[31] = 64'b1111111111111111111111111111111100000000000000000000000000000000;
	  assign write_buffer[32] = 64'b1111111111111111111111111111111110000000000000000000000000000000;
	  assign write_buffer[33] = 64'b1111111111111111111111111111111111000000000000000000000000000000;
	  assign write_buffer[34] = 64'b1111111111111111111111111111111111100000000000000000000000000000;
	  assign write_buffer[35] = 64'b1111111111111111111111111111111111110000000000000000000000000000;
	  assign write_buffer[36] = 64'b1111111111111111111111111111111111111000000000000000000000000000;
	  assign write_buffer[37] = 64'b1111111111111111111111111111111111111100000000000000000000000000;
	  assign write_buffer[38] = 64'b1111111111111111111111111111111111111110000000000000000000000000;
	  assign write_buffer[39] = 64'b1111111111111111111111111111111111111111000000000000000000000000;
	  assign write_buffer[40] = 64'b1111111111111111111111111111111111111111100000000000000000000000;
	  assign write_buffer[41] = 64'b1111111111111111111111111111111111111111110000000000000000000000;
	  assign write_buffer[42] = 64'b1111111111111111111111111111111111111111111000000000000000000000;
	  assign write_buffer[43] = 64'b1111111111111111111111111111111111111111111100000000000000000000;
	  assign write_buffer[44] = 64'b1111111111111111111111111111111111111111111110000000000000000000;
	  assign write_buffer[45] = 64'b1111111111111111111111111111111111111111111111000000000000000000;
	  assign write_buffer[46] = 64'b1111111111111111111111111111111111111111111111100000000000000000;
	  assign write_buffer[47] = 64'b1111111111111111111111111111111111111111111111110000000000000000;
	  assign write_buffer[48] = 64'b1111111111111111111111111111111111111111111111111000000000000000;
	  assign write_buffer[49] = 64'b1111111111111111111111111111111111111111111111111100000000000000;
	  assign write_buffer[50] = 64'b1111111111111111111111111111111111111111111111111110000000000000;
	  assign write_buffer[51] = 64'b1111111111111111111111111111111111111111111111111111000000000000;
	  assign write_buffer[52] = 64'b1111111111111111111111111111111111111111111111111111100000000000;
	  assign write_buffer[53] = 64'b1111111111111111111111111111111111111111111111111111110000000000;
	  assign write_buffer[54] = 64'b1111111111111111111111111111111111111111111111111111111000000000;
	  assign write_buffer[55] = 64'b1111111111111111111111111111111111111111111111111111111100000000;
	  assign write_buffer[56] = 64'b1111111111111111111111111111111111111111111111111111111110000000;
	  assign write_buffer[57] = 64'b1111111111111111111111111111111111111111111111111111111111000000;
	  assign write_buffer[58] = 64'b1111111111111111111111111111111111111111111111111111111111100000;
	  assign write_buffer[59] = 64'b1111111111111111111111111111111111111111111111111111111111110000;
	  assign write_buffer[60] = 64'b1111111111111111111111111111111111111111111111111111111111111000;
	  assign write_buffer[61] = 64'b1111111111111111111111111111111111111111111111111111111111111100;
	  assign write_buffer[62] = 64'b1111111111111111111111111111111111111111111111111111111111111110;
	  assign write_buffer[63] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 
	 
	  logic [63:0] row_0_in;
	  logic [63:0] row_1_in;
	

	  logic [5:0] row_0_sel;
	  logic [5:0] row_1_sel;
	  assign row_0_sel = addr;
	  assign row_1_sel = addr+32;
	  
	  logic read_en;

	  DisplayController #(.WIDTH(WIDTH)) DisplayControllerTest(clk, reset, row_0_in, row_1_in, addr, OE, latch, r0_out, r1_out, g0_out, g1_out, b0_out, b1_out,sck,read_en);
	 


	  TESTMEMReadControl  TestMem(clk,reset,read_en,row_0_sel,row_1_sel,write_buffer, row_0_in,row_1_in );
endmodule



//////////////////////////////////////////////////////////////////////
//							TESTEBRDisplay	MODULE					//
//							A TESTING MODULE						//
//////////////////////////////////////////////////////////////////////
module TESTMemoryDisplay #(WIDTH=4)   (input logic clk,
									input logic reset,
									output logic r0_out,
									output logic r1_out,
									output logic g0_out,
									output logic g1_out,
									output logic b0_out,
									output logic b1_out,  
									output logic latch,
									output logic OE,
									output logic sck,
									output logic [4:0] addr);
	
	logic [5:0] data_count;
	logic  [5:0] data_frame [63:0];
	logic data_ready;
	
	//data_count counter
	always_ff @(posedge clk)begin
		if(reset) data_count = 0;
		else data_count = data_count+1;
	end
	
	//stuff for "simulating" SPI in hardware
	always_ff @(posedge clk)begin
		if(data_count==4  )begin
			data_ready <= 1;
			for(int i = 0; i<64;i=i+1)begin
				data_frame[i] <= i+data_count;
			end
		end
		else data_ready <= 0;
	end
	
	MemoryDisplay #(.WIDTH(WIDTH)) TestMod(clk, reset, data_frame, data_ready, r0_out, r1_out, g0_out, g1_out, b0_out, b1_out, latch, OE, sck, addr);
	
endmodule




module TESTMEMReadControl  (input logic clk,
						input logic reset,
						input logic r_en,
						input logic [5:0] row_0_sel,
						input logic [5:0] row_1_sel,
						input logic [63:0] write_buffer [63:0], 
						output logic [63:0] row_0,
						output logic [63:0]row_1 );
	logic [63:0] read_buffer [63:0];
	always_ff @(posedge clk) begin
		if(r_en)begin
			row_0 <= read_buffer[row_0_sel];
			row_1 <= read_buffer[row_1_sel];
		end
		read_buffer<=write_buffer;
	end	
endmodule

